module sigmoid (
    input clk,
    input [11:0] x,
    output [11:0] score
);
    always @ (posedge clk) begin
        

endmodule