module notgate(a,b);
    input a;
    output b;

    assign b = ~a;
endmodule